* Extracted by KLayout with SG13G2 LVS runset on : 12/05/2025 15:47

.SUBCKT 2NmosSch
X$1 \$1 Vdd G1 Vout power_switch_nmos
X$2 \$1 GND G2 Vout power_switch_nmos
.ENDS 2NmosSch

.SUBCKT power_switch_nmos \$1 \$2 \$3 \$14
X$1 \$1 \$2 power_switch_nmos_isolbox
X$2 \$1 \$2 power_switch_nmos_gr3
X$3 \$2 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3
+ \$3 \$3 \$3 \$3 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14
+ \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14
+ \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14
+ \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 power_switch_nmos_side
X$4 \$2 \$3 power_switch_nmos_gate_trunk
X$5 \$2 power_switch_nmos_gr1
X$6 \$2 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3 \$3
+ \$3 \$3 \$3 \$3 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14
+ \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14
+ \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14
+ \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 \$14 power_switch_nmos_side
.ENDS power_switch_nmos

.SUBCKT power_switch_nmos_gr3 \$1 \$2
.ENDS power_switch_nmos_gr3

.SUBCKT power_switch_nmos_isolbox \$1 \$5
.ENDS power_switch_nmos_isolbox

.SUBCKT power_switch_nmos_gr1 \$1
.ENDS power_switch_nmos_gr1

.SUBCKT power_switch_nmos_gate_trunk \$1 \$2
.ENDS power_switch_nmos_gate_trunk

.SUBCKT power_switch_nmos_side \$1 \$2 \$3 \$4 \$5 \$6 \$7 \$8 \$9 \$10 \$11
+ \$12 \$13 \$14 \$15 \$16 \$17 \$18 \$19 \$20 \$21 \$I698 \$I688 \$I659 \$I640
+ \$I621 \$I602 \$I583 \$I564 \$I545 \$I526 \$I507 \$I488 \$I469 \$I450 \$I431
+ \$I412 \$I393 \$I374 \$I355 \$I336 \$I317 \$I298 \$I279 \$I260 \$I241 \$I222
+ \$I203 \$I192 \$I165 \$I164 \$I163 \$I162 \$I161 \$I160 \$I159 \$I158 \$I157
+ \$I156 \$I155 \$I154 \$I153 \$I152 \$I151 \$I150 \$I149 \$I148 \$I147 \$I146
+ \$I145 \$I144 \$I143 \$I142 \$I141 \$I132
X$1 \$1 \$19 \$21 \$I132 \$I203 \$I222 \$I241 \$I260 \$I279 \$I298 \$I317
+ \$I336 \$I355 \$I374 \$I393 \$I412 \$I431 \$I450 \$I469 \$I488 \$I507 \$I526
+ \$I545 \$I564 \$I583 \$I602 \$I621 \$I640 \$I659 power_switch_nblock
X$2 \$1 \$18 \$20 \$I192 \$I165 \$I164 \$I163 \$I162 \$I161 \$I160 \$I159
+ \$I158 \$I157 \$I156 \$I155 \$I154 \$I153 \$I152 \$I151 \$I150 \$I149 \$I148
+ \$I147 \$I146 \$I145 \$I144 \$I143 \$I142 \$I141 power_switch_nblock
X$3 \$1 \$I141 \$1 via_m4m5_long$1
X$4 \$1 \$I142 \$1 via_m4m5_long$1
X$5 \$1 \$I143 \$1 via_m4m5_long$1
X$6 \$1 \$I144 \$1 via_m4m5_long$1
X$7 \$1 \$I145 \$1 via_m4m5_long$1
X$8 \$1 \$I146 \$1 via_m4m5_long$1
X$9 \$1 \$I147 \$1 via_m4m5_long$1
X$10 \$1 \$I148 \$1 via_m4m5_long$1
X$11 \$1 \$I149 \$1 via_m4m5_long$1
X$12 \$1 \$I150 \$1 via_m4m5_long$1
X$13 \$1 \$I151 \$1 via_m4m5_long$1
X$14 \$1 \$I152 \$1 via_m4m5_long$1
X$15 \$1 \$I153 \$1 via_m4m5_long$1
X$16 \$1 \$I154 \$1 via_m4m5_long$1
X$17 \$1 \$I155 \$1 via_m4m5_long$1
X$18 \$1 \$I156 \$1 via_m4m5_long$1
X$19 \$1 \$I157 \$1 via_m4m5_long$1
X$20 \$1 \$I158 \$1 via_m4m5_long$1
X$21 \$1 \$I159 \$1 via_m4m5_long$1
X$22 \$1 \$I160 \$1 via_m4m5_long$1
X$23 \$1 \$I161 \$1 via_m4m5_long$1
X$24 \$1 \$I162 \$1 via_m4m5_long$1
X$25 \$1 \$I163 \$1 via_m4m5_long$1
X$26 \$1 \$I164 \$1 via_m4m5_long$1
X$27 \$1 \$I165 \$1 via_m4m5_long$1
X$28 \$1 \$I192 \$1 via_m4m5_long$1
X$29 \$1 \$16 \$18 \$I192 \$I165 \$I164 \$I163 \$I162 \$I161 \$I160 \$I159
+ \$I158 \$I157 \$I156 \$I155 \$I154 \$I153 \$I152 \$I151 \$I150 \$I149 \$I148
+ \$I147 \$I146 \$I145 \$I144 \$I143 \$I142 \$I141 power_switch_nblock
X$30 \$1 \$17 \$19 \$I132 \$I203 \$I222 \$I241 \$I260 \$I279 \$I298 \$I317
+ \$I336 \$I355 \$I374 \$I393 \$I412 \$I431 \$I450 \$I469 \$I488 \$I507 \$I526
+ \$I545 \$I564 \$I583 \$I602 \$I621 \$I640 \$I659 power_switch_nblock
X$31 \$1 \$14 \$16 \$I192 \$I165 \$I164 \$I163 \$I162 \$I161 \$I160 \$I159
+ \$I158 \$I157 \$I156 \$I155 \$I154 \$I153 \$I152 \$I151 \$I150 \$I149 \$I148
+ \$I147 \$I146 \$I145 \$I144 \$I143 \$I142 \$I141 power_switch_nblock
X$32 \$1 \$15 \$17 \$I132 \$I203 \$I222 \$I241 \$I260 \$I279 \$I298 \$I317
+ \$I336 \$I355 \$I374 \$I393 \$I412 \$I431 \$I450 \$I469 \$I488 \$I507 \$I526
+ \$I545 \$I564 \$I583 \$I602 \$I621 \$I640 \$I659 power_switch_nblock
X$33 \$1 \$12 \$14 \$I192 \$I165 \$I164 \$I163 \$I162 \$I161 \$I160 \$I159
+ \$I158 \$I157 \$I156 \$I155 \$I154 \$I153 \$I152 \$I151 \$I150 \$I149 \$I148
+ \$I147 \$I146 \$I145 \$I144 \$I143 \$I142 \$I141 power_switch_nblock
X$34 \$1 \$13 \$15 \$I132 \$I203 \$I222 \$I241 \$I260 \$I279 \$I298 \$I317
+ \$I336 \$I355 \$I374 \$I393 \$I412 \$I431 \$I450 \$I469 \$I488 \$I507 \$I526
+ \$I545 \$I564 \$I583 \$I602 \$I621 \$I640 \$I659 power_switch_nblock
X$35 \$1 \$10 \$12 \$I192 \$I165 \$I164 \$I163 \$I162 \$I161 \$I160 \$I159
+ \$I158 \$I157 \$I156 \$I155 \$I154 \$I153 \$I152 \$I151 \$I150 \$I149 \$I148
+ \$I147 \$I146 \$I145 \$I144 \$I143 \$I142 \$I141 power_switch_nblock
X$36 \$1 \$11 \$13 \$I132 \$I203 \$I222 \$I241 \$I260 \$I279 \$I298 \$I317
+ \$I336 \$I355 \$I374 \$I393 \$I412 \$I431 \$I450 \$I469 \$I488 \$I507 \$I526
+ \$I545 \$I564 \$I583 \$I602 \$I621 \$I640 \$I659 power_switch_nblock
X$37 \$1 \$8 \$10 \$I192 \$I165 \$I164 \$I163 \$I162 \$I161 \$I160 \$I159
+ \$I158 \$I157 \$I156 \$I155 \$I154 \$I153 \$I152 \$I151 \$I150 \$I149 \$I148
+ \$I147 \$I146 \$I145 \$I144 \$I143 \$I142 \$I141 power_switch_nblock
X$38 \$1 \$9 \$11 \$I132 \$I203 \$I222 \$I241 \$I260 \$I279 \$I298 \$I317
+ \$I336 \$I355 \$I374 \$I393 \$I412 \$I431 \$I450 \$I469 \$I488 \$I507 \$I526
+ \$I545 \$I564 \$I583 \$I602 \$I621 \$I640 \$I659 power_switch_nblock
X$39 \$1 \$6 \$8 \$I192 \$I165 \$I164 \$I163 \$I162 \$I161 \$I160 \$I159 \$I158
+ \$I157 \$I156 \$I155 \$I154 \$I153 \$I152 \$I151 \$I150 \$I149 \$I148 \$I147
+ \$I146 \$I145 \$I144 \$I143 \$I142 \$I141 power_switch_nblock
X$40 \$1 \$7 \$9 \$I132 \$I203 \$I222 \$I241 \$I260 \$I279 \$I298 \$I317 \$I336
+ \$I355 \$I374 \$I393 \$I412 \$I431 \$I450 \$I469 \$I488 \$I507 \$I526 \$I545
+ \$I564 \$I583 \$I602 \$I621 \$I640 \$I659 power_switch_nblock
X$41 \$1 \$4 \$6 \$I192 \$I165 \$I164 \$I163 \$I162 \$I161 \$I160 \$I159 \$I158
+ \$I157 \$I156 \$I155 \$I154 \$I153 \$I152 \$I151 \$I150 \$I149 \$I148 \$I147
+ \$I146 \$I145 \$I144 \$I143 \$I142 \$I141 power_switch_nblock
X$42 \$1 \$5 \$7 \$I132 \$I203 \$I222 \$I241 \$I260 \$I279 \$I298 \$I317 \$I336
+ \$I355 \$I374 \$I393 \$I412 \$I431 \$I450 \$I469 \$I488 \$I507 \$I526 \$I545
+ \$I564 \$I583 \$I602 \$I621 \$I640 \$I659 power_switch_nblock
X$43 \$1 \$2 \$4 \$I192 \$I165 \$I164 \$I163 \$I162 \$I161 \$I160 \$I159 \$I158
+ \$I157 \$I156 \$I155 \$I154 \$I153 \$I152 \$I151 \$I150 \$I149 \$I148 \$I147
+ \$I146 \$I145 \$I144 \$I143 \$I142 \$I141 power_switch_nblock
X$44 \$1 \$3 \$5 \$I132 \$I203 \$I222 \$I241 \$I260 \$I279 \$I298 \$I317 \$I336
+ \$I355 \$I374 \$I393 \$I412 \$I431 \$I450 \$I469 \$I488 \$I507 \$I526 \$I545
+ \$I564 \$I583 \$I602 \$I621 \$I640 \$I659 power_switch_nblock
X$45 \$1 \$I698 \$2 \$I192 \$I165 \$I164 \$I163 \$I162 \$I161 \$I160 \$I159
+ \$I158 \$I157 \$I156 \$I155 \$I154 \$I153 \$I152 \$I151 \$I150 \$I149 \$I148
+ \$I147 \$I146 \$I145 \$I144 \$I143 \$I142 \$I141 power_switch_nblock
X$46 \$1 \$I688 \$3 \$I132 \$I203 \$I222 \$I241 \$I260 \$I279 \$I298 \$I317
+ \$I336 \$I355 \$I374 \$I393 \$I412 \$I431 \$I450 \$I469 \$I488 \$I507 \$I526
+ \$I545 \$I564 \$I583 \$I602 \$I621 \$I640 \$I659 power_switch_nblock
X$47 \$1 \$I659 \$1 via_m4m5_long$1
X$48 \$1 \$I640 \$1 via_m4m5_long$1
X$49 \$1 \$I621 \$1 via_m4m5_long$1
X$50 \$1 \$I602 \$1 via_m4m5_long$1
X$51 \$1 \$I583 \$1 via_m4m5_long$1
X$52 \$1 \$I564 \$1 via_m4m5_long$1
X$53 \$1 \$I545 \$1 via_m4m5_long$1
X$54 \$1 \$I526 \$1 via_m4m5_long$1
X$55 \$1 \$I507 \$1 via_m4m5_long$1
X$56 \$1 \$I488 \$1 via_m4m5_long$1
X$57 \$1 \$I469 \$1 via_m4m5_long$1
X$58 \$1 \$I450 \$1 via_m4m5_long$1
X$59 \$1 \$I431 \$1 via_m4m5_long$1
X$60 \$1 \$I412 \$1 via_m4m5_long$1
X$61 \$1 \$I393 \$1 via_m4m5_long$1
X$62 \$1 \$I374 \$1 via_m4m5_long$1
X$63 \$1 \$I355 \$1 via_m4m5_long$1
X$64 \$1 \$I336 \$1 via_m4m5_long$1
X$65 \$1 \$I317 \$1 via_m4m5_long$1
X$66 \$1 \$I298 \$1 via_m4m5_long$1
X$67 \$1 \$I279 \$1 via_m4m5_long$1
X$68 \$1 \$I260 \$1 via_m4m5_long$1
X$69 \$1 \$I241 \$1 via_m4m5_long$1
X$70 \$1 \$I222 \$1 via_m4m5_long$1
X$71 \$1 \$I203 \$1 via_m4m5_long$1
X$72 \$1 \$I132 \$1 via_m4m5_long$1
.ENDS power_switch_nmos_side

.SUBCKT via_m4m5_long$1 \$1 \$2 \$3
.ENDS via_m4m5_long$1

.SUBCKT power_switch_nblock \$1 \$I133 \$I132 \$I56 \$I55 \$I54 \$I53 \$I52
+ \$I51 \$I50 \$I49 \$I48 \$I47 \$I46 \$I45 \$I44 \$I43 \$I42 \$I41 \$I40 \$I39
+ \$I38 \$I37 \$I36 \$I35 \$I34 \$I33 \$I32 \$I31
X$1 \$I133 \$1 \$I56 \$1 \$I55 \$1 \$I54 \$1 \$I53 \$1 \$I52 \$1 \$I51 \$1
+ \$I50 \$1 \$I49 \$1 \$I48 \$1 \$I47 \$1 \$I46 \$1 \$I45 \$1 \$I44 \$1 \$I43
+ \$1 \$I42 \$1 \$I41 \$1 \$I40 \$1 \$I39 \$1 \$I38 \$1 \$I37 \$1 \$I36 \$1
+ \$I35 \$1 \$I34 \$1 \$I33 \$1 \$I32 \$1 \$I31 \$1 power_switch_nfingers
X$2 \$1 \$1 \$I56 via_m3m4_1x2
X$3 \$I132 \$I31 \$1 \$I32 \$1 \$I33 \$1 \$I34 \$1 \$I35 \$1 \$I36 \$1 \$I37
+ \$1 \$I38 \$1 \$I39 \$1 \$I40 \$1 \$I41 \$1 \$I42 \$1 \$I43 \$1 \$I44 \$1
+ \$I45 \$1 \$I46 \$1 \$I47 \$1 \$I48 \$1 \$I49 \$1 \$I50 \$1 \$I51 \$1 \$I52
+ \$1 \$I53 \$1 \$I54 \$1 \$I55 \$1 \$I56 \$1 \$1 power_switch_nfingers
X$4 \$1 Unnamed_45933b9e
X$5 \$1 \$1 \$I31 via_m3m4_1x2
X$6 \$1 \$1 \$I32 via_m3m4_1x2
X$7 \$1 \$1 \$I33 via_m3m4_1x2
X$8 \$1 \$1 \$I34 via_m3m4_1x2
X$9 \$1 \$1 \$I35 via_m3m4_1x2
X$10 \$1 \$1 \$I36 via_m3m4_1x2
X$11 \$1 \$1 \$I37 via_m3m4_1x2
X$12 \$1 \$1 \$I38 via_m3m4_1x2
X$13 \$1 \$1 \$I39 via_m3m4_1x2
X$14 \$1 \$1 \$I40 via_m3m4_1x2
X$15 \$1 \$1 \$I41 via_m3m4_1x2
X$16 \$1 \$1 \$I42 via_m3m4_1x2
X$17 \$1 \$1 \$I43 via_m3m4_1x2
X$18 \$1 \$1 \$I44 via_m3m4_1x2
X$19 \$1 \$1 \$I45 via_m3m4_1x2
X$20 \$1 \$1 \$I46 via_m3m4_1x2
X$21 \$1 \$1 \$I47 via_m3m4_1x2
X$22 \$1 \$1 \$I48 via_m3m4_1x2
X$23 \$1 \$1 \$I49 via_m3m4_1x2
X$24 \$1 \$1 \$I50 via_m3m4_1x2
X$25 \$1 \$1 \$I51 via_m3m4_1x2
X$26 \$1 \$1 \$I52 via_m3m4_1x2
X$27 \$1 \$1 \$I53 via_m3m4_1x2
X$28 \$1 \$1 \$I54 via_m3m4_1x2
X$29 \$1 \$1 \$I55 via_m3m4_1x2
.ENDS power_switch_nblock

.SUBCKT via_m3m4_1x2 \$1 \$2 \$3
.ENDS via_m3m4_1x2

.SUBCKT Unnamed_45933b9e \$1
.ENDS Unnamed_45933b9e

.SUBCKT power_switch_nfingers \$1 \$2 \$3 \$4 \$5 \$6 \$7 \$8 \$9 \$10 \$11
+ \$12 \$13 \$14 \$15 \$16 \$17 \$18 \$19 \$20 \$21 \$22 \$23 \$24 \$25 \$26
+ \$27 \$28 \$29 \$30 \$31 \$32 \$33 \$34 \$35 \$36 \$37 \$38 \$39 \$40 \$41
+ \$42 \$43 \$44 \$45 \$46 \$47 \$48 \$49 \$50 \$51 \$52 \$53 \$54
X$1 \$2 \$54 via_array_cda5390a
X$2 \$3 \$54 via_array_cda5390a
X$3 \$4 \$54 via_array_cda5390a
X$4 \$5 \$54 via_array_cda5390a
X$5 \$6 \$54 via_array_cda5390a
X$6 \$7 \$54 via_array_cda5390a
X$7 \$8 \$54 via_array_cda5390a
X$8 \$9 \$54 via_array_cda5390a
X$9 \$10 \$54 via_array_cda5390a
X$10 \$11 \$54 via_array_cda5390a
X$11 \$12 \$54 via_array_cda5390a
X$12 \$13 \$54 via_array_cda5390a
X$13 \$14 \$54 via_array_cda5390a
X$14 \$15 \$54 via_array_cda5390a
X$15 \$16 \$54 via_array_cda5390a
X$16 \$17 \$54 via_array_cda5390a
X$17 \$18 \$54 via_array_cda5390a
X$18 \$19 \$54 via_array_cda5390a
X$19 \$20 \$54 via_array_cda5390a
X$20 \$21 \$54 via_array_cda5390a
X$21 \$22 \$54 via_array_cda5390a
X$22 \$23 \$54 via_array_cda5390a
X$23 \$24 \$54 via_array_cda5390a
X$24 \$25 \$54 via_array_cda5390a
X$25 \$26 \$54 via_array_cda5390a
X$26 \$27 \$54 via_array_cda5390a
X$27 \$28 \$54 via_array_cda5390a
X$28 \$29 \$54 via_array_cda5390a
X$29 \$30 \$54 via_array_cda5390a
X$30 \$31 \$54 via_array_cda5390a
X$31 \$32 \$54 via_array_cda5390a
X$32 \$33 \$54 via_array_cda5390a
X$33 \$34 \$54 via_array_cda5390a
X$34 \$35 \$54 via_array_cda5390a
X$35 \$36 \$54 via_array_cda5390a
X$36 \$37 \$54 via_array_cda5390a
X$37 \$38 \$54 via_array_cda5390a
X$38 \$39 \$54 via_array_cda5390a
X$39 \$40 \$54 via_array_cda5390a
X$40 \$41 \$54 via_array_cda5390a
X$41 \$42 \$54 via_array_cda5390a
X$42 \$43 \$54 via_array_cda5390a
X$43 \$44 \$54 via_array_cda5390a
X$44 \$45 \$54 via_array_cda5390a
X$45 \$46 \$54 via_array_cda5390a
X$46 \$47 \$54 via_array_cda5390a
X$47 \$48 \$54 via_array_cda5390a
X$48 \$49 \$54 via_array_cda5390a
X$49 \$50 \$54 via_array_cda5390a
X$50 \$51 \$54 via_array_cda5390a
X$51 \$52 \$54 via_array_cda5390a
X$52 \$53 \$54 via_array_cda5390a
M$1 \$2 \$1 \$3 \$54 sg13_hv_nmos L=0.45u W=10u AS=7.7p AD=3.5p PS=21.54u
+ PD=10.7u
M$2 \$3 \$1 \$4 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$3 \$4 \$1 \$5 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$4 \$5 \$1 \$6 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$5 \$6 \$1 \$7 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$6 \$7 \$1 \$8 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$7 \$8 \$1 \$9 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$8 \$9 \$1 \$10 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$9 \$10 \$1 \$11 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$10 \$11 \$1 \$12 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$11 \$12 \$1 \$13 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$12 \$13 \$1 \$14 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$13 \$14 \$1 \$15 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$14 \$15 \$1 \$16 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$15 \$16 \$1 \$17 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$16 \$17 \$1 \$18 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$17 \$18 \$1 \$19 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$18 \$19 \$1 \$20 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$19 \$20 \$1 \$21 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$20 \$21 \$1 \$22 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$21 \$22 \$1 \$23 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$22 \$23 \$1 \$24 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$23 \$24 \$1 \$25 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$24 \$25 \$1 \$26 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$25 \$26 \$1 \$27 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$26 \$27 \$1 \$28 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$27 \$28 \$1 \$29 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$28 \$29 \$1 \$30 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$29 \$30 \$1 \$31 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$30 \$31 \$1 \$32 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$31 \$32 \$1 \$33 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$32 \$33 \$1 \$34 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$33 \$34 \$1 \$35 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$34 \$35 \$1 \$36 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$35 \$36 \$1 \$37 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$36 \$37 \$1 \$38 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$37 \$38 \$1 \$39 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$38 \$39 \$1 \$40 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$39 \$40 \$1 \$41 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$40 \$41 \$1 \$42 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$41 \$42 \$1 \$43 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$42 \$43 \$1 \$44 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$43 \$44 \$1 \$45 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$44 \$45 \$1 \$46 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$45 \$46 \$1 \$47 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$46 \$47 \$1 \$48 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$47 \$48 \$1 \$49 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$48 \$49 \$1 \$50 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$49 \$50 \$1 \$51 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$50 \$51 \$1 \$52 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=3.5p PS=10.7u
+ PD=10.7u
M$51 \$52 \$1 \$53 \$54 sg13_hv_nmos L=0.45u W=10u AS=3.5p AD=7.7p PS=10.7u
+ PD=21.54u
.ENDS power_switch_nfingers

.SUBCKT via_array_cda5390a \$1 \$2
.ENDS via_array_cda5390a
